library ieee;
use ieee.std_logic_1164.all;

package mac_package is
		constant W : integer := 8;
end; -- mac package
