library ieee;
use ieee.std_logic_1164.all;

package bram_package is
		constant W	:	integer := 32;
		constant L	:	integer :=1024;
end; -- blockram package
