Library ieee;
Use ieee.std_logic_1164.all;
Entity or2 is
Port (
	A : in std_logic;
	B : in std_logic;
	Z : out std_logic
);
end or2;
architecture dataflow of or2 is
begin
Z <= A or B;
end dataflow;
